module IDU(

);
endmodule
