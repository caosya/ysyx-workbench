module ALU(

);
endmodule
