module Reg(

);
endmodule
