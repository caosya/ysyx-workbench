module Mem(

);
endmodule
